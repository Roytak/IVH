--------------------------------------------------------------------------------
-- IVH Project
-- Author: Roman Janota
-- Date : 08/05/2022
--	File : anewspaper_pack.vhd
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package newspaper_pack is

type DIRECTION_T is (DIR_LEFT,DIR_RIGHT,DIR_ANIM);

end newspaper_pack;

package body newspaper_pack is

end newspaper_pack;
